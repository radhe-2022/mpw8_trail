magic
tech sky130A
magscale 1 2
timestamp 1672346171
<< nwell >>
rect 1066 77509 78882 77830
rect 1066 76421 78882 76987
rect 1066 75333 78882 75899
rect 1066 74245 78882 74811
rect 1066 73157 78882 73723
rect 1066 72069 78882 72635
rect 1066 70981 78882 71547
rect 1066 69893 78882 70459
rect 1066 68805 78882 69371
rect 1066 67717 78882 68283
rect 1066 66629 78882 67195
rect 1066 65541 78882 66107
rect 1066 64453 78882 65019
rect 1066 63365 78882 63931
rect 1066 62277 78882 62843
rect 1066 61189 78882 61755
rect 1066 60101 78882 60667
rect 1066 59013 78882 59579
rect 1066 57925 78882 58491
rect 1066 56837 78882 57403
rect 1066 55749 78882 56315
rect 1066 54661 78882 55227
rect 1066 53573 78882 54139
rect 1066 52485 78882 53051
rect 1066 51397 78882 51963
rect 1066 50309 78882 50875
rect 1066 49221 78882 49787
rect 1066 48133 78882 48699
rect 1066 47045 78882 47611
rect 1066 45957 78882 46523
rect 1066 44869 78882 45435
rect 1066 43781 78882 44347
rect 1066 42693 78882 43259
rect 1066 41605 78882 42171
rect 1066 40517 78882 41083
rect 1066 39429 78882 39995
rect 1066 38341 78882 38907
rect 1066 37253 78882 37819
rect 1066 36165 78882 36731
rect 1066 35077 78882 35643
rect 1066 33989 78882 34555
rect 1066 32901 78882 33467
rect 1066 31813 78882 32379
rect 1066 30725 78882 31291
rect 1066 29637 78882 30203
rect 1066 28549 78882 29115
rect 1066 27461 78882 28027
rect 1066 26373 78882 26939
rect 1066 25285 78882 25851
rect 1066 24197 78882 24763
rect 1066 23109 78882 23675
rect 1066 22021 78882 22587
rect 1066 20933 78882 21499
rect 1066 19845 78882 20411
rect 1066 18757 78882 19323
rect 1066 17669 78882 18235
rect 1066 16581 78882 17147
rect 1066 15493 78882 16059
rect 1066 14405 78882 14971
rect 1066 13317 78882 13883
rect 1066 12229 78882 12795
rect 1066 11141 78882 11707
rect 1066 10053 78882 10619
rect 1066 8965 78882 9531
rect 1066 7877 78882 8443
rect 1066 6789 78882 7355
rect 1066 5701 78882 6267
rect 1066 4613 78882 5179
rect 1066 3525 78882 4091
rect 1066 2437 78882 3003
<< obsli1 >>
rect 1104 2159 78844 77809
<< obsm1 >>
rect 1104 2048 78844 77840
<< metal2 >>
rect 5170 79200 5226 80000
rect 15106 79200 15162 80000
rect 25042 79200 25098 80000
rect 34978 79200 35034 80000
rect 44914 79200 44970 80000
rect 54850 79200 54906 80000
rect 64786 79200 64842 80000
rect 74722 79200 74778 80000
rect 2410 0 2466 800
rect 5538 0 5594 800
rect 8666 0 8722 800
rect 11794 0 11850 800
rect 14922 0 14978 800
rect 18050 0 18106 800
rect 21178 0 21234 800
rect 24306 0 24362 800
rect 27434 0 27490 800
rect 30562 0 30618 800
rect 33690 0 33746 800
rect 36818 0 36874 800
rect 39946 0 40002 800
rect 43074 0 43130 800
rect 46202 0 46258 800
rect 49330 0 49386 800
rect 52458 0 52514 800
rect 55586 0 55642 800
rect 58714 0 58770 800
rect 61842 0 61898 800
rect 64970 0 65026 800
rect 68098 0 68154 800
rect 71226 0 71282 800
rect 74354 0 74410 800
rect 77482 0 77538 800
<< obsm2 >>
rect 2412 79144 5114 79200
rect 5282 79144 15050 79200
rect 15218 79144 24986 79200
rect 25154 79144 34922 79200
rect 35090 79144 44858 79200
rect 45026 79144 54794 79200
rect 54962 79144 64730 79200
rect 64898 79144 74666 79200
rect 74834 79144 77536 79200
rect 2412 856 77536 79144
rect 2522 800 5482 856
rect 5650 800 8610 856
rect 8778 800 11738 856
rect 11906 800 14866 856
rect 15034 800 17994 856
rect 18162 800 21122 856
rect 21290 800 24250 856
rect 24418 800 27378 856
rect 27546 800 30506 856
rect 30674 800 33634 856
rect 33802 800 36762 856
rect 36930 800 39890 856
rect 40058 800 43018 856
rect 43186 800 46146 856
rect 46314 800 49274 856
rect 49442 800 52402 856
rect 52570 800 55530 856
rect 55698 800 58658 856
rect 58826 800 61786 856
rect 61954 800 64914 856
rect 65082 800 68042 856
rect 68210 800 71170 856
rect 71338 800 74298 856
rect 74466 800 77426 856
<< obsm3 >>
rect 2773 2143 77083 77825
<< metal4 >>
rect 4208 2128 4528 77840
rect 19568 2128 19888 77840
rect 34928 2128 35248 77840
rect 50288 2128 50608 77840
rect 65648 2128 65968 77840
<< obsm4 >>
rect 13307 3435 19488 77485
rect 19968 3435 34848 77485
rect 35328 3435 50208 77485
rect 50688 3435 61949 77485
<< labels >>
rlabel metal2 s 25042 79200 25098 80000 6 clk
port 1 nsew signal input
rlabel metal2 s 15106 79200 15162 80000 6 execute
port 2 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 input_val[0]
port 3 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 input_val[1]
port 4 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 input_val[2]
port 5 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 input_val[3]
port 6 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 input_val[4]
port 7 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 input_val[5]
port 8 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 input_val[6]
port 9 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 input_val[7]
port 10 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 out[0]
port 11 nsew signal output
rlabel metal2 s 58714 0 58770 800 6 out[10]
port 12 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 out[11]
port 13 nsew signal output
rlabel metal2 s 64970 0 65026 800 6 out[12]
port 14 nsew signal output
rlabel metal2 s 68098 0 68154 800 6 out[13]
port 15 nsew signal output
rlabel metal2 s 71226 0 71282 800 6 out[14]
port 16 nsew signal output
rlabel metal2 s 74354 0 74410 800 6 out[15]
port 17 nsew signal output
rlabel metal2 s 77482 0 77538 800 6 out[16]
port 18 nsew signal output
rlabel metal2 s 30562 0 30618 800 6 out[1]
port 19 nsew signal output
rlabel metal2 s 33690 0 33746 800 6 out[2]
port 20 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 out[3]
port 21 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 out[4]
port 22 nsew signal output
rlabel metal2 s 43074 0 43130 800 6 out[5]
port 23 nsew signal output
rlabel metal2 s 46202 0 46258 800 6 out[6]
port 24 nsew signal output
rlabel metal2 s 49330 0 49386 800 6 out[7]
port 25 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 out[8]
port 26 nsew signal output
rlabel metal2 s 55586 0 55642 800 6 out[9]
port 27 nsew signal output
rlabel metal2 s 5170 79200 5226 80000 6 reset
port 28 nsew signal input
rlabel metal2 s 34978 79200 35034 80000 6 sel_in[0]
port 29 nsew signal input
rlabel metal2 s 44914 79200 44970 80000 6 sel_in[1]
port 30 nsew signal input
rlabel metal2 s 54850 79200 54906 80000 6 sel_in[2]
port 31 nsew signal input
rlabel metal2 s 64786 79200 64842 80000 6 sel_out[0]
port 32 nsew signal input
rlabel metal2 s 74722 79200 74778 80000 6 sel_out[1]
port 33 nsew signal input
rlabel metal4 s 4208 2128 4528 77840 6 vccd1
port 34 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 77840 6 vccd1
port 34 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 77840 6 vccd1
port 34 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 77840 6 vssd1
port 35 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 77840 6 vssd1
port 35 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 80000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 11979850
string GDS_FILE /home/radhe/project/mpw8_trail/openlane/matrix_multiply/runs/22_12_30_01_54/results/signoff/matrix_multiply.magic.gds
string GDS_START 809888
<< end >>

